`timescale 1ns / 1ps
/////////////////////
module dff(d,clk,q);
output reg q;
input d,clk;
always@(posedge clk)
begin
q<=d;
end

endmodule
